module normalizeFrac(num, a, b);
input[23:0] a;
input[4:0] num;
output reg[23:0] b;
always @(a or num)
begin
case(num)	
	5'b00000: b={a[23:0]};
	5'b00001: b={a[22:0],1'b0};
	5'b00010: b={a[21:0],2'b0};
	5'b00011: b={a[20:0],3'b0};
	5'b00100: b={a[19:0],4'b0};
	5'b00101: b={a[18:0],5'b0};
	5'b00110: b={a[17:0],6'b0};
	5'b00111: b={a[16:0],7'b0};
	5'b01000: b={a[15:0],8'b0};
	5'b01001: b={a[14:0],9'b0};
	5'b01010: b={a[13:0],10'b0};
	5'b01011: b={a[12:0],11'b0};
	5'b01100: b={a[11:0],12'b0};
	5'b01101: b={a[10:0],13'b0};
	5'b01110: b={a[9:0],14'b0};
	5'b01111: b={a[8:0],15'b0};
	5'b10000: b={a[7:0],16'b0};
	5'b10001: b={a[6:0],17'b0};
	5'b10010: b={a[5:0],18'b0};
	5'b10011: b={a[4:0],19'b0};
	5'b10100: b={a[3:0],20'b0};
	5'b10101: b={a[2:0],21'b0};
	5'b10110: b={a[1:0],22'b0};
	5'b10111: b={a[0],23'b0};
	default: b=24'b0;
endcase
end
endmodule