module fadder(x, y, cin, s, cout);
input x, y, cin;
output s, cout;
wire m1,m2,m3;
xor(m1,x,y);
xor(s,cin,m1);
and(m2,cin,m1);
and(m3,x,y);
or(cout,m3,m2);
endmodule

module mux2(a1, b1, s1, f1);   
input a1, b1, s1;
output f1;
wire m4,m5,m6;
	not(m4,s1);
	and(m5,m4,a1);
	and(m6,s1,b1);
	or(f1,m5,m6);
endmodule

module add_csa(a,b,ci,s,co);
	input wire [24:0]a,b;
	input wire ci;
	output wire [24:0]s;
	output wire co;
	wire [24:0] temp0,temp1,c0,c1,t;
	xor(t[0], b[0], ci);
	xor(t[1], b[1], ci);
	xor(t[2], b[2], ci);
	xor(t[3], b[3], ci);
	xor(t[4], b[4], ci);
	xor(t[5], b[5], ci); 
	xor(t[6], b[6], ci);
	xor(t[7], b[7], ci);
	xor(t[8], b[8], ci);
	xor(t[9], b[9], ci);
	xor(t[10], b[10], ci);
	xor(t[11], b[11], ci);
	xor(t[12], b[12], ci);
	xor(t[13], b[13], ci); 
	xor(t[14], b[14], ci);
	xor(t[15], b[15], ci);
	xor(t[16], b[16], ci);
	xor(t[17], b[17], ci);
	xor(t[18], b[18], ci);
	xor(t[19], b[19], ci);
	xor(t[20], b[20], ci);
	xor(t[21], b[21], ci); 
	xor(t[22], b[22], ci);
	xor(t[23], b[23], ci);
	xor(t[24], b[24], ci);
//carry 0
	fadder fa000(a[0] ,t[0] ,1'b0  ,temp0[0] ,c0[0] );
	fadder fa001(a[1] ,t[1] ,c0[0] ,temp0[1] ,c0[1] );	
	fadder fa002(a[2] ,t[2] ,c0[1] ,temp0[2] ,c0[2] );	
	fadder fa003(a[3] ,t[3] ,c0[2] ,temp0[3] ,c0[3] );
	fadder fa004(a[4] ,t[4] ,c0[3] ,temp0[4] ,c0[4] );	
	fadder fa005(a[5] ,t[5] ,c0[4] ,temp0[5] ,c0[5] );	
	fadder fa006(a[6] ,t[6] ,c0[5] ,temp0[6] ,c0[6] );
	fadder fa007(a[7] ,t[7] ,c0[6] ,temp0[7] ,c0[7] );
	fadder fa008(a[8] ,t[8] ,c0[7] ,temp0[8] ,c0[8] );	
	fadder fa009(a[9] ,t[9] ,c0[8] ,temp0[9] ,c0[9] );	
	fadder fa010(a[10],t[10],c0[9] ,temp0[10],c0[10]);
	fadder fa011(a[11],t[11],c0[10],temp0[11],c0[11]);	
	fadder fa012(a[12],t[12],c0[11],temp0[12],c0[12]);	
	fadder fa013(a[13],t[13],c0[12],temp0[13],c0[13]);
	fadder fa014(a[14],t[14],c0[13],temp0[14],c0[14]);
	fadder fa015(a[15],t[15],c0[14],temp0[15],c0[15]);	
	fadder fa016(a[16],t[16],c0[15],temp0[16],c0[16]);	
	fadder fa017(a[17],t[17],c0[16],temp0[17],c0[17]);
	fadder fa018(a[18],t[18],c0[17],temp0[18],c0[18]);	
	fadder fa019(a[19],t[19],c0[18],temp0[19],c0[19]);	
	fadder fa020(a[20],t[20],c0[19],temp0[20],c0[20]);
	fadder fa021(a[21],t[21],c0[20],temp0[21],c0[21]);
	fadder fa022(a[22],t[22],c0[21],temp0[22],c0[22]);
	fadder fa023(a[23],t[23],c0[22],temp0[23],c0[23]);
	fadder fa024(a[24],t[24],c0[23],temp0[24],c0[24]);

//carry 1
	fadder fa100(a[0] ,t[0] ,1'b1  ,temp1[0] ,c1[0] );
	fadder fa101(a[1] ,t[1] ,c1[0] ,temp1[1] ,c1[1] );	
	fadder fa102(a[2] ,t[2] ,c1[1] ,temp1[2] ,c1[2] );	
	fadder fa103(a[3] ,t[3] ,c1[2] ,temp1[3] ,c1[3] );
	fadder fa104(a[4] ,t[4] ,c1[3] ,temp1[4] ,c1[4] );	
	fadder fa105(a[5] ,t[5] ,c1[4] ,temp1[5] ,c1[5] );	
	fadder fa106(a[6] ,t[6] ,c1[5] ,temp1[6] ,c1[6] );
	fadder fa107(a[7] ,t[7] ,c1[6] ,temp1[7] ,c1[7] );
	fadder fa108(a[8] ,t[8] ,c1[7] ,temp1[8] ,c1[8] );	
	fadder fa109(a[9] ,t[9] ,c1[8] ,temp1[9] ,c1[9] );	
	fadder fa110(a[10],t[10],c1[9] ,temp1[10],c1[10]);
	fadder fa111(a[11],t[11],c1[10],temp1[11],c1[11]);	
	fadder fa112(a[12],t[12],c1[11],temp1[12],c1[12]);	
	fadder fa113(a[13],t[13],c1[12],temp1[13],c1[13]);
	fadder fa114(a[14],t[14],c1[13],temp1[14],c1[14]);
	fadder fa115(a[15],t[15],c1[14],temp1[15],c1[15]);	
	fadder fa116(a[16],t[16],c1[15],temp1[16],c1[16]);	
	fadder fa117(a[17],t[17],c1[16],temp1[17],c1[17]);
	fadder fa118(a[18],t[18],c1[17],temp1[18],c1[18]);	
	fadder fa119(a[19],t[19],c1[18],temp1[19],c1[19]);	
	fadder fa120(a[20],t[20],c1[19],temp1[20],c1[20]);
	fadder fa121(a[21],t[21],c1[20],temp1[21],c1[21]);
	fadder fa122(a[22],t[22],c1[21],temp1[22],c1[22]);
	fadder fa123(a[23],t[23],c1[22],temp1[23],c1[23]);
	fadder fa124(a[24],t[24],c1[23],temp1[24],c1[24]);
//mux carry
	mux2 mux_c(c0[23],c1[23],ci,co);
//mux sum
	mux2 muxs0 (temp0[0] ,temp1[0] ,ci,s[0] );
	mux2 muxs1 (temp0[1] ,temp1[1] ,ci,s[1] );	
	mux2 muxs2 (temp0[2] ,temp1[2] ,ci,s[2] );	
	mux2 muxs3 (temp0[3] ,temp1[3] ,ci,s[3] );
	mux2 muxs4 (temp0[4] ,temp1[4] ,ci,s[4] );
	mux2 muxs5 (temp0[5] ,temp1[5] ,ci,s[5] );	
	mux2 muxs6 (temp0[6] ,temp1[6] ,ci,s[6] );	
	mux2 muxs7 (temp0[7] ,temp1[7] ,ci,s[7] );
	mux2 muxs8 (temp0[8] ,temp1[8] ,ci,s[8] );
	mux2 muxs9 (temp0[9] ,temp1[9] ,ci,s[9] );	
	mux2 muxs10(temp0[10],temp1[10],ci,s[10]);	
	mux2 muxs11(temp0[11],temp1[11],ci,s[11]);
	mux2 muxs12(temp0[12],temp1[12],ci,s[12]);
	mux2 muxs13(temp0[13],temp1[13],ci,s[13]);	
	mux2 muxs14(temp0[14],temp1[14],ci,s[14]);	
	mux2 muxs15(temp0[15],temp1[15],ci,s[15]);
	mux2 muxs16(temp0[16],temp1[16],ci,s[16]);
	mux2 muxs17(temp0[17],temp1[17],ci,s[17]);	
	mux2 muxs18(temp0[18],temp1[18],ci,s[18]);	
	mux2 muxs19(temp0[19],temp1[19],ci,s[19]);
	mux2 muxs20(temp0[20],temp1[20],ci,s[20]);
	mux2 muxs21(temp0[21],temp1[21],ci,s[21]);	
	mux2 muxs22(temp0[22],temp1[22],ci,s[22]);	
	mux2 muxs23(temp0[23],temp1[23],ci,s[23]);	
	mux2 muxs24(temp0[24],temp1[24],ci,s[24]);
endmodule
