module main(a,b,sel,s);
input[31:0] a,b;
input sel;
output[31:0] s;
wire[7:0] exo;
wire siga, sigb;
wire[2:0] ctro;
wire alhb, cout2;
wire[7:0] numshift;
wire[23:0] shiftrout, swapoa, swapob;
wire[22:0] muxo1, muxo2; 
wire[24:0] signialu, neg2out;
wire[23:0] normalin,normalfracout;
wire[4:0] normalo;
SmallAlu Smallalu1(a[30:23],b[30:23],numshift,alhb);
control controlu(alhb,ctro);
mux2_23b mux23_1(a[22:0],b[22:0],ctro[1],muxo1);
mux2_23b mux23_2(a[22:0],b[22:0],ctro[0],muxo2);
mux2_8b mux2_1(a[30:23],b[30:23],ctro[2],exo);
Shiftright Dichphai(numshift,{1'b1,muxo1},shiftrout);
Swap_ab Swap1(shiftrout,{1'b1,muxo2},alhb,swapoa,swapob);
Bigalu alusignificant(swapoa,swapob,sel,signialu,cout2);
bu2ifam bu2ifneg(signialu,neg2out);
normalize detectbit1(neg2out[24:1],normalo);
normalizeFrac normalfrac1(normalo,neg2out[24:1],normalfracout);
normalizeExpo normalexpo1(normalo,exo,s[30:23]);
assign s[22:0]=normalfracout[22:0];
Xacdinhdau Dau1(s[31],sel,cout2,a[31],b[31]);
endmodule