library verilog;
use verilog.vl_types.all;
entity check0 is
    port(
        a               : in     vl_logic_vector(7 downto 0);
        f               : out    vl_logic
    );
end check0;
